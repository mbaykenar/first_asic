magic
tech sky130A
magscale 1 2
timestamp 1658211152
<< obsli1 >>
rect 1104 2159 198812 197489
<< obsm1 >>
rect 14 2128 199718 197520
<< metal2 >>
rect 18 199200 74 200000
rect 3238 199200 3294 200000
rect 7102 199200 7158 200000
rect 10322 199200 10378 200000
rect 13542 199200 13598 200000
rect 16762 199200 16818 200000
rect 19982 199200 20038 200000
rect 23202 199200 23258 200000
rect 26422 199200 26478 200000
rect 29642 199200 29698 200000
rect 32862 199200 32918 200000
rect 36082 199200 36138 200000
rect 39302 199200 39358 200000
rect 42522 199200 42578 200000
rect 46386 199200 46442 200000
rect 49606 199200 49662 200000
rect 52826 199200 52882 200000
rect 56046 199200 56102 200000
rect 59266 199200 59322 200000
rect 62486 199200 62542 200000
rect 65706 199200 65762 200000
rect 68926 199200 68982 200000
rect 72146 199200 72202 200000
rect 75366 199200 75422 200000
rect 78586 199200 78642 200000
rect 81806 199200 81862 200000
rect 85670 199200 85726 200000
rect 88890 199200 88946 200000
rect 92110 199200 92166 200000
rect 95330 199200 95386 200000
rect 98550 199200 98606 200000
rect 101770 199200 101826 200000
rect 104990 199200 105046 200000
rect 108210 199200 108266 200000
rect 111430 199200 111486 200000
rect 114650 199200 114706 200000
rect 117870 199200 117926 200000
rect 121090 199200 121146 200000
rect 124954 199200 125010 200000
rect 128174 199200 128230 200000
rect 131394 199200 131450 200000
rect 134614 199200 134670 200000
rect 137834 199200 137890 200000
rect 141054 199200 141110 200000
rect 144274 199200 144330 200000
rect 147494 199200 147550 200000
rect 150714 199200 150770 200000
rect 153934 199200 153990 200000
rect 157154 199200 157210 200000
rect 160374 199200 160430 200000
rect 164238 199200 164294 200000
rect 167458 199200 167514 200000
rect 170678 199200 170734 200000
rect 173898 199200 173954 200000
rect 177118 199200 177174 200000
rect 180338 199200 180394 200000
rect 183558 199200 183614 200000
rect 186778 199200 186834 200000
rect 189998 199200 190054 200000
rect 193218 199200 193274 200000
rect 196438 199200 196494 200000
rect 199658 199200 199714 200000
rect 18 0 74 800
rect 3238 0 3294 800
rect 6458 0 6514 800
rect 9678 0 9734 800
rect 12898 0 12954 800
rect 16118 0 16174 800
rect 19338 0 19394 800
rect 22558 0 22614 800
rect 25778 0 25834 800
rect 28998 0 29054 800
rect 32218 0 32274 800
rect 35438 0 35494 800
rect 39302 0 39358 800
rect 42522 0 42578 800
rect 45742 0 45798 800
rect 48962 0 49018 800
rect 52182 0 52238 800
rect 55402 0 55458 800
rect 58622 0 58678 800
rect 61842 0 61898 800
rect 65062 0 65118 800
rect 68282 0 68338 800
rect 71502 0 71558 800
rect 74722 0 74778 800
rect 78586 0 78642 800
rect 81806 0 81862 800
rect 85026 0 85082 800
rect 88246 0 88302 800
rect 91466 0 91522 800
rect 94686 0 94742 800
rect 97906 0 97962 800
rect 101126 0 101182 800
rect 104346 0 104402 800
rect 107566 0 107622 800
rect 110786 0 110842 800
rect 114006 0 114062 800
rect 117870 0 117926 800
rect 121090 0 121146 800
rect 124310 0 124366 800
rect 127530 0 127586 800
rect 130750 0 130806 800
rect 133970 0 134026 800
rect 137190 0 137246 800
rect 140410 0 140466 800
rect 143630 0 143686 800
rect 146850 0 146906 800
rect 150070 0 150126 800
rect 153290 0 153346 800
rect 157154 0 157210 800
rect 160374 0 160430 800
rect 163594 0 163650 800
rect 166814 0 166870 800
rect 170034 0 170090 800
rect 173254 0 173310 800
rect 176474 0 176530 800
rect 179694 0 179750 800
rect 182914 0 182970 800
rect 186134 0 186190 800
rect 189354 0 189410 800
rect 192574 0 192630 800
rect 196438 0 196494 800
rect 199658 0 199714 800
<< obsm2 >>
rect 130 199144 3182 199322
rect 3350 199144 7046 199322
rect 7214 199144 10266 199322
rect 10434 199144 13486 199322
rect 13654 199144 16706 199322
rect 16874 199144 19926 199322
rect 20094 199144 23146 199322
rect 23314 199144 26366 199322
rect 26534 199144 29586 199322
rect 29754 199144 32806 199322
rect 32974 199144 36026 199322
rect 36194 199144 39246 199322
rect 39414 199144 42466 199322
rect 42634 199144 46330 199322
rect 46498 199144 49550 199322
rect 49718 199144 52770 199322
rect 52938 199144 55990 199322
rect 56158 199144 59210 199322
rect 59378 199144 62430 199322
rect 62598 199144 65650 199322
rect 65818 199144 68870 199322
rect 69038 199144 72090 199322
rect 72258 199144 75310 199322
rect 75478 199144 78530 199322
rect 78698 199144 81750 199322
rect 81918 199144 85614 199322
rect 85782 199144 88834 199322
rect 89002 199144 92054 199322
rect 92222 199144 95274 199322
rect 95442 199144 98494 199322
rect 98662 199144 101714 199322
rect 101882 199144 104934 199322
rect 105102 199144 108154 199322
rect 108322 199144 111374 199322
rect 111542 199144 114594 199322
rect 114762 199144 117814 199322
rect 117982 199144 121034 199322
rect 121202 199144 124898 199322
rect 125066 199144 128118 199322
rect 128286 199144 131338 199322
rect 131506 199144 134558 199322
rect 134726 199144 137778 199322
rect 137946 199144 140998 199322
rect 141166 199144 144218 199322
rect 144386 199144 147438 199322
rect 147606 199144 150658 199322
rect 150826 199144 153878 199322
rect 154046 199144 157098 199322
rect 157266 199144 160318 199322
rect 160486 199144 164182 199322
rect 164350 199144 167402 199322
rect 167570 199144 170622 199322
rect 170790 199144 173842 199322
rect 174010 199144 177062 199322
rect 177230 199144 180282 199322
rect 180450 199144 183502 199322
rect 183670 199144 186722 199322
rect 186890 199144 189942 199322
rect 190110 199144 193162 199322
rect 193330 199144 196382 199322
rect 196550 199144 199602 199322
rect 20 856 199712 199144
rect 130 734 3182 856
rect 3350 734 6402 856
rect 6570 734 9622 856
rect 9790 734 12842 856
rect 13010 734 16062 856
rect 16230 734 19282 856
rect 19450 734 22502 856
rect 22670 734 25722 856
rect 25890 734 28942 856
rect 29110 734 32162 856
rect 32330 734 35382 856
rect 35550 734 39246 856
rect 39414 734 42466 856
rect 42634 734 45686 856
rect 45854 734 48906 856
rect 49074 734 52126 856
rect 52294 734 55346 856
rect 55514 734 58566 856
rect 58734 734 61786 856
rect 61954 734 65006 856
rect 65174 734 68226 856
rect 68394 734 71446 856
rect 71614 734 74666 856
rect 74834 734 78530 856
rect 78698 734 81750 856
rect 81918 734 84970 856
rect 85138 734 88190 856
rect 88358 734 91410 856
rect 91578 734 94630 856
rect 94798 734 97850 856
rect 98018 734 101070 856
rect 101238 734 104290 856
rect 104458 734 107510 856
rect 107678 734 110730 856
rect 110898 734 113950 856
rect 114118 734 117814 856
rect 117982 734 121034 856
rect 121202 734 124254 856
rect 124422 734 127474 856
rect 127642 734 130694 856
rect 130862 734 133914 856
rect 134082 734 137134 856
rect 137302 734 140354 856
rect 140522 734 143574 856
rect 143742 734 146794 856
rect 146962 734 150014 856
rect 150182 734 153234 856
rect 153402 734 157098 856
rect 157266 734 160318 856
rect 160486 734 163538 856
rect 163706 734 166758 856
rect 166926 734 169978 856
rect 170146 734 173198 856
rect 173366 734 176418 856
rect 176586 734 179638 856
rect 179806 734 182858 856
rect 183026 734 186078 856
rect 186246 734 189298 856
rect 189466 734 192518 856
rect 192686 734 196382 856
rect 196550 734 199602 856
<< metal3 >>
rect 0 196528 800 196648
rect 199200 195848 200000 195968
rect 0 193128 800 193248
rect 199200 192448 200000 192568
rect 0 189728 800 189848
rect 199200 189048 200000 189168
rect 0 186328 800 186448
rect 199200 185648 200000 185768
rect 0 182928 800 183048
rect 199200 182248 200000 182368
rect 0 179528 800 179648
rect 199200 178848 200000 178968
rect 0 176128 800 176248
rect 199200 175448 200000 175568
rect 0 172728 800 172848
rect 199200 172048 200000 172168
rect 0 169328 800 169448
rect 199200 168648 200000 168768
rect 0 165928 800 166048
rect 199200 165248 200000 165368
rect 0 161848 800 161968
rect 199200 161848 200000 161968
rect 0 158448 800 158568
rect 199200 157768 200000 157888
rect 0 155048 800 155168
rect 199200 154368 200000 154488
rect 0 151648 800 151768
rect 199200 150968 200000 151088
rect 0 148248 800 148368
rect 199200 147568 200000 147688
rect 0 144848 800 144968
rect 199200 144168 200000 144288
rect 0 141448 800 141568
rect 199200 140768 200000 140888
rect 0 138048 800 138168
rect 199200 137368 200000 137488
rect 0 134648 800 134768
rect 199200 133968 200000 134088
rect 0 131248 800 131368
rect 199200 130568 200000 130688
rect 0 127848 800 127968
rect 199200 127168 200000 127288
rect 0 124448 800 124568
rect 199200 123768 200000 123888
rect 0 120368 800 120488
rect 199200 120368 200000 120488
rect 0 116968 800 117088
rect 199200 116288 200000 116408
rect 0 113568 800 113688
rect 199200 112888 200000 113008
rect 0 110168 800 110288
rect 199200 109488 200000 109608
rect 0 106768 800 106888
rect 199200 106088 200000 106208
rect 0 103368 800 103488
rect 199200 102688 200000 102808
rect 0 99968 800 100088
rect 199200 99288 200000 99408
rect 0 96568 800 96688
rect 199200 95888 200000 96008
rect 0 93168 800 93288
rect 199200 92488 200000 92608
rect 0 89768 800 89888
rect 199200 89088 200000 89208
rect 0 86368 800 86488
rect 199200 85688 200000 85808
rect 0 82968 800 83088
rect 199200 82288 200000 82408
rect 0 78888 800 79008
rect 199200 78888 200000 79008
rect 0 75488 800 75608
rect 199200 74808 200000 74928
rect 0 72088 800 72208
rect 199200 71408 200000 71528
rect 0 68688 800 68808
rect 199200 68008 200000 68128
rect 0 65288 800 65408
rect 199200 64608 200000 64728
rect 0 61888 800 62008
rect 199200 61208 200000 61328
rect 0 58488 800 58608
rect 199200 57808 200000 57928
rect 0 55088 800 55208
rect 199200 54408 200000 54528
rect 0 51688 800 51808
rect 199200 51008 200000 51128
rect 0 48288 800 48408
rect 199200 47608 200000 47728
rect 0 44888 800 45008
rect 199200 44208 200000 44328
rect 0 41488 800 41608
rect 199200 40808 200000 40928
rect 0 37408 800 37528
rect 199200 37408 200000 37528
rect 0 34008 800 34128
rect 199200 33328 200000 33448
rect 0 30608 800 30728
rect 199200 29928 200000 30048
rect 0 27208 800 27328
rect 199200 26528 200000 26648
rect 0 23808 800 23928
rect 199200 23128 200000 23248
rect 0 20408 800 20528
rect 199200 19728 200000 19848
rect 0 17008 800 17128
rect 199200 16328 200000 16448
rect 0 13608 800 13728
rect 199200 12928 200000 13048
rect 0 10208 800 10328
rect 199200 9528 200000 9648
rect 0 6808 800 6928
rect 199200 6128 200000 6248
rect 0 3408 800 3528
rect 199200 2728 200000 2848
<< obsm3 >>
rect 800 196728 199200 197505
rect 880 196448 199200 196728
rect 800 196048 199200 196448
rect 800 195768 199120 196048
rect 800 193328 199200 195768
rect 880 193048 199200 193328
rect 800 192648 199200 193048
rect 800 192368 199120 192648
rect 800 189928 199200 192368
rect 880 189648 199200 189928
rect 800 189248 199200 189648
rect 800 188968 199120 189248
rect 800 186528 199200 188968
rect 880 186248 199200 186528
rect 800 185848 199200 186248
rect 800 185568 199120 185848
rect 800 183128 199200 185568
rect 880 182848 199200 183128
rect 800 182448 199200 182848
rect 800 182168 199120 182448
rect 800 179728 199200 182168
rect 880 179448 199200 179728
rect 800 179048 199200 179448
rect 800 178768 199120 179048
rect 800 176328 199200 178768
rect 880 176048 199200 176328
rect 800 175648 199200 176048
rect 800 175368 199120 175648
rect 800 172928 199200 175368
rect 880 172648 199200 172928
rect 800 172248 199200 172648
rect 800 171968 199120 172248
rect 800 169528 199200 171968
rect 880 169248 199200 169528
rect 800 168848 199200 169248
rect 800 168568 199120 168848
rect 800 166128 199200 168568
rect 880 165848 199200 166128
rect 800 165448 199200 165848
rect 800 165168 199120 165448
rect 800 162048 199200 165168
rect 880 161768 199120 162048
rect 800 158648 199200 161768
rect 880 158368 199200 158648
rect 800 157968 199200 158368
rect 800 157688 199120 157968
rect 800 155248 199200 157688
rect 880 154968 199200 155248
rect 800 154568 199200 154968
rect 800 154288 199120 154568
rect 800 151848 199200 154288
rect 880 151568 199200 151848
rect 800 151168 199200 151568
rect 800 150888 199120 151168
rect 800 148448 199200 150888
rect 880 148168 199200 148448
rect 800 147768 199200 148168
rect 800 147488 199120 147768
rect 800 145048 199200 147488
rect 880 144768 199200 145048
rect 800 144368 199200 144768
rect 800 144088 199120 144368
rect 800 141648 199200 144088
rect 880 141368 199200 141648
rect 800 140968 199200 141368
rect 800 140688 199120 140968
rect 800 138248 199200 140688
rect 880 137968 199200 138248
rect 800 137568 199200 137968
rect 800 137288 199120 137568
rect 800 134848 199200 137288
rect 880 134568 199200 134848
rect 800 134168 199200 134568
rect 800 133888 199120 134168
rect 800 131448 199200 133888
rect 880 131168 199200 131448
rect 800 130768 199200 131168
rect 800 130488 199120 130768
rect 800 128048 199200 130488
rect 880 127768 199200 128048
rect 800 127368 199200 127768
rect 800 127088 199120 127368
rect 800 124648 199200 127088
rect 880 124368 199200 124648
rect 800 123968 199200 124368
rect 800 123688 199120 123968
rect 800 120568 199200 123688
rect 880 120288 199120 120568
rect 800 117168 199200 120288
rect 880 116888 199200 117168
rect 800 116488 199200 116888
rect 800 116208 199120 116488
rect 800 113768 199200 116208
rect 880 113488 199200 113768
rect 800 113088 199200 113488
rect 800 112808 199120 113088
rect 800 110368 199200 112808
rect 880 110088 199200 110368
rect 800 109688 199200 110088
rect 800 109408 199120 109688
rect 800 106968 199200 109408
rect 880 106688 199200 106968
rect 800 106288 199200 106688
rect 800 106008 199120 106288
rect 800 103568 199200 106008
rect 880 103288 199200 103568
rect 800 102888 199200 103288
rect 800 102608 199120 102888
rect 800 100168 199200 102608
rect 880 99888 199200 100168
rect 800 99488 199200 99888
rect 800 99208 199120 99488
rect 800 96768 199200 99208
rect 880 96488 199200 96768
rect 800 96088 199200 96488
rect 800 95808 199120 96088
rect 800 93368 199200 95808
rect 880 93088 199200 93368
rect 800 92688 199200 93088
rect 800 92408 199120 92688
rect 800 89968 199200 92408
rect 880 89688 199200 89968
rect 800 89288 199200 89688
rect 800 89008 199120 89288
rect 800 86568 199200 89008
rect 880 86288 199200 86568
rect 800 85888 199200 86288
rect 800 85608 199120 85888
rect 800 83168 199200 85608
rect 880 82888 199200 83168
rect 800 82488 199200 82888
rect 800 82208 199120 82488
rect 800 79088 199200 82208
rect 880 78808 199120 79088
rect 800 75688 199200 78808
rect 880 75408 199200 75688
rect 800 75008 199200 75408
rect 800 74728 199120 75008
rect 800 72288 199200 74728
rect 880 72008 199200 72288
rect 800 71608 199200 72008
rect 800 71328 199120 71608
rect 800 68888 199200 71328
rect 880 68608 199200 68888
rect 800 68208 199200 68608
rect 800 67928 199120 68208
rect 800 65488 199200 67928
rect 880 65208 199200 65488
rect 800 64808 199200 65208
rect 800 64528 199120 64808
rect 800 62088 199200 64528
rect 880 61808 199200 62088
rect 800 61408 199200 61808
rect 800 61128 199120 61408
rect 800 58688 199200 61128
rect 880 58408 199200 58688
rect 800 58008 199200 58408
rect 800 57728 199120 58008
rect 800 55288 199200 57728
rect 880 55008 199200 55288
rect 800 54608 199200 55008
rect 800 54328 199120 54608
rect 800 51888 199200 54328
rect 880 51608 199200 51888
rect 800 51208 199200 51608
rect 800 50928 199120 51208
rect 800 48488 199200 50928
rect 880 48208 199200 48488
rect 800 47808 199200 48208
rect 800 47528 199120 47808
rect 800 45088 199200 47528
rect 880 44808 199200 45088
rect 800 44408 199200 44808
rect 800 44128 199120 44408
rect 800 41688 199200 44128
rect 880 41408 199200 41688
rect 800 41008 199200 41408
rect 800 40728 199120 41008
rect 800 37608 199200 40728
rect 880 37328 199120 37608
rect 800 34208 199200 37328
rect 880 33928 199200 34208
rect 800 33528 199200 33928
rect 800 33248 199120 33528
rect 800 30808 199200 33248
rect 880 30528 199200 30808
rect 800 30128 199200 30528
rect 800 29848 199120 30128
rect 800 27408 199200 29848
rect 880 27128 199200 27408
rect 800 26728 199200 27128
rect 800 26448 199120 26728
rect 800 24008 199200 26448
rect 880 23728 199200 24008
rect 800 23328 199200 23728
rect 800 23048 199120 23328
rect 800 20608 199200 23048
rect 880 20328 199200 20608
rect 800 19928 199200 20328
rect 800 19648 199120 19928
rect 800 17208 199200 19648
rect 880 16928 199200 17208
rect 800 16528 199200 16928
rect 800 16248 199120 16528
rect 800 13808 199200 16248
rect 880 13528 199200 13808
rect 800 13128 199200 13528
rect 800 12848 199120 13128
rect 800 10408 199200 12848
rect 880 10128 199200 10408
rect 800 9728 199200 10128
rect 800 9448 199120 9728
rect 800 7008 199200 9448
rect 880 6728 199200 7008
rect 800 6328 199200 6728
rect 800 6048 199120 6328
rect 800 3608 199200 6048
rect 880 3328 199200 3608
rect 800 2928 199200 3328
rect 800 2648 199120 2928
rect 800 2143 199200 2648
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
rect 111728 2128 112048 197520
rect 127088 2128 127408 197520
rect 142448 2128 142768 197520
rect 157808 2128 158128 197520
rect 173168 2128 173488 197520
rect 188528 2128 188848 197520
<< obsm4 >>
rect 64827 2483 65568 197165
rect 66048 2483 80928 197165
rect 81408 2483 96288 197165
rect 96768 2483 111648 197165
rect 112128 2483 118805 197165
<< metal5 >>
rect 1104 189114 198812 189434
rect 1104 173796 198812 174116
rect 1104 158478 198812 158798
rect 1104 143160 198812 143480
rect 1104 127842 198812 128162
rect 1104 112524 198812 112844
rect 1104 97206 198812 97526
rect 1104 81888 198812 82208
rect 1104 66570 198812 66890
rect 1104 51252 198812 51572
rect 1104 35934 198812 36254
rect 1104 20616 198812 20936
rect 1104 5298 198812 5618
<< labels >>
rlabel metal2 s 160374 0 160430 800 6 alu_adder_ext_i[0]
port 1 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 alu_adder_ext_i[10]
port 2 nsew signal input
rlabel metal3 s 199200 182248 200000 182368 6 alu_adder_ext_i[11]
port 3 nsew signal input
rlabel metal3 s 199200 71408 200000 71528 6 alu_adder_ext_i[12]
port 4 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 alu_adder_ext_i[13]
port 5 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 alu_adder_ext_i[14]
port 6 nsew signal input
rlabel metal2 s 134614 199200 134670 200000 6 alu_adder_ext_i[15]
port 7 nsew signal input
rlabel metal2 s 68926 199200 68982 200000 6 alu_adder_ext_i[16]
port 8 nsew signal input
rlabel metal2 s 170678 199200 170734 200000 6 alu_adder_ext_i[17]
port 9 nsew signal input
rlabel metal2 s 18 199200 74 200000 6 alu_adder_ext_i[18]
port 10 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 alu_adder_ext_i[19]
port 11 nsew signal input
rlabel metal3 s 199200 61208 200000 61328 6 alu_adder_ext_i[1]
port 12 nsew signal input
rlabel metal3 s 0 193128 800 193248 6 alu_adder_ext_i[20]
port 13 nsew signal input
rlabel metal2 s 42522 199200 42578 200000 6 alu_adder_ext_i[21]
port 14 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 alu_adder_ext_i[22]
port 15 nsew signal input
rlabel metal2 s 36082 199200 36138 200000 6 alu_adder_ext_i[23]
port 16 nsew signal input
rlabel metal3 s 199200 102688 200000 102808 6 alu_adder_ext_i[24]
port 17 nsew signal input
rlabel metal3 s 199200 165248 200000 165368 6 alu_adder_ext_i[25]
port 18 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 alu_adder_ext_i[26]
port 19 nsew signal input
rlabel metal2 s 59266 199200 59322 200000 6 alu_adder_ext_i[27]
port 20 nsew signal input
rlabel metal2 s 78586 199200 78642 200000 6 alu_adder_ext_i[28]
port 21 nsew signal input
rlabel metal2 s 164238 199200 164294 200000 6 alu_adder_ext_i[29]
port 22 nsew signal input
rlabel metal2 s 98550 199200 98606 200000 6 alu_adder_ext_i[2]
port 23 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 alu_adder_ext_i[30]
port 24 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 alu_adder_ext_i[31]
port 25 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 alu_adder_ext_i[32]
port 26 nsew signal input
rlabel metal3 s 199200 82288 200000 82408 6 alu_adder_ext_i[33]
port 27 nsew signal input
rlabel metal2 s 186134 0 186190 800 6 alu_adder_ext_i[3]
port 28 nsew signal input
rlabel metal3 s 0 155048 800 155168 6 alu_adder_ext_i[4]
port 29 nsew signal input
rlabel metal3 s 199200 178848 200000 178968 6 alu_adder_ext_i[5]
port 30 nsew signal input
rlabel metal3 s 199200 26528 200000 26648 6 alu_adder_ext_i[6]
port 31 nsew signal input
rlabel metal2 s 150714 199200 150770 200000 6 alu_adder_ext_i[7]
port 32 nsew signal input
rlabel metal3 s 199200 92488 200000 92608 6 alu_adder_ext_i[8]
port 33 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 alu_adder_ext_i[9]
port 34 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 alu_adder_i[0]
port 35 nsew signal input
rlabel metal2 s 32862 199200 32918 200000 6 alu_adder_i[10]
port 36 nsew signal input
rlabel metal2 s 121090 199200 121146 200000 6 alu_adder_i[11]
port 37 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 alu_adder_i[12]
port 38 nsew signal input
rlabel metal3 s 199200 137368 200000 137488 6 alu_adder_i[13]
port 39 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 alu_adder_i[14]
port 40 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 alu_adder_i[15]
port 41 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 alu_adder_i[16]
port 42 nsew signal input
rlabel metal2 s 183558 199200 183614 200000 6 alu_adder_i[17]
port 43 nsew signal input
rlabel metal3 s 199200 99288 200000 99408 6 alu_adder_i[18]
port 44 nsew signal input
rlabel metal3 s 0 138048 800 138168 6 alu_adder_i[19]
port 45 nsew signal input
rlabel metal3 s 199200 40808 200000 40928 6 alu_adder_i[1]
port 46 nsew signal input
rlabel metal3 s 199200 106088 200000 106208 6 alu_adder_i[20]
port 47 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 alu_adder_i[21]
port 48 nsew signal input
rlabel metal2 s 49606 199200 49662 200000 6 alu_adder_i[22]
port 49 nsew signal input
rlabel metal2 s 131394 199200 131450 200000 6 alu_adder_i[23]
port 50 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 alu_adder_i[24]
port 51 nsew signal input
rlabel metal3 s 199200 68008 200000 68128 6 alu_adder_i[25]
port 52 nsew signal input
rlabel metal2 s 13542 199200 13598 200000 6 alu_adder_i[26]
port 53 nsew signal input
rlabel metal3 s 199200 130568 200000 130688 6 alu_adder_i[27]
port 54 nsew signal input
rlabel metal3 s 0 169328 800 169448 6 alu_adder_i[28]
port 55 nsew signal input
rlabel metal2 s 111430 199200 111486 200000 6 alu_adder_i[29]
port 56 nsew signal input
rlabel metal2 s 117870 199200 117926 200000 6 alu_adder_i[2]
port 57 nsew signal input
rlabel metal2 s 19982 199200 20038 200000 6 alu_adder_i[30]
port 58 nsew signal input
rlabel metal2 s 85670 199200 85726 200000 6 alu_adder_i[31]
port 59 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 alu_adder_i[3]
port 60 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 alu_adder_i[4]
port 61 nsew signal input
rlabel metal2 s 179694 0 179750 800 6 alu_adder_i[5]
port 62 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 alu_adder_i[6]
port 63 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 alu_adder_i[7]
port 64 nsew signal input
rlabel metal3 s 199200 120368 200000 120488 6 alu_adder_i[8]
port 65 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 alu_adder_i[9]
port 66 nsew signal input
rlabel metal3 s 0 165928 800 166048 6 alu_operand_a_o[0]
port 67 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 alu_operand_a_o[10]
port 68 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 alu_operand_a_o[11]
port 69 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 alu_operand_a_o[12]
port 70 nsew signal output
rlabel metal2 s 92110 199200 92166 200000 6 alu_operand_a_o[13]
port 71 nsew signal output
rlabel metal2 s 95330 199200 95386 200000 6 alu_operand_a_o[14]
port 72 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 alu_operand_a_o[15]
port 73 nsew signal output
rlabel metal2 s 186778 199200 186834 200000 6 alu_operand_a_o[16]
port 74 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 alu_operand_a_o[17]
port 75 nsew signal output
rlabel metal2 s 153290 0 153346 800 6 alu_operand_a_o[18]
port 76 nsew signal output
rlabel metal3 s 199200 12928 200000 13048 6 alu_operand_a_o[19]
port 77 nsew signal output
rlabel metal3 s 199200 19728 200000 19848 6 alu_operand_a_o[1]
port 78 nsew signal output
rlabel metal3 s 199200 37408 200000 37528 6 alu_operand_a_o[20]
port 79 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 alu_operand_a_o[21]
port 80 nsew signal output
rlabel metal2 s 157154 199200 157210 200000 6 alu_operand_a_o[22]
port 81 nsew signal output
rlabel metal3 s 199200 154368 200000 154488 6 alu_operand_a_o[23]
port 82 nsew signal output
rlabel metal3 s 199200 51008 200000 51128 6 alu_operand_a_o[24]
port 83 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 alu_operand_a_o[25]
port 84 nsew signal output
rlabel metal2 s 166814 0 166870 800 6 alu_operand_a_o[26]
port 85 nsew signal output
rlabel metal2 s 72146 199200 72202 200000 6 alu_operand_a_o[27]
port 86 nsew signal output
rlabel metal3 s 199200 23128 200000 23248 6 alu_operand_a_o[28]
port 87 nsew signal output
rlabel metal2 s 189998 199200 190054 200000 6 alu_operand_a_o[29]
port 88 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 alu_operand_a_o[2]
port 89 nsew signal output
rlabel metal3 s 199200 6128 200000 6248 6 alu_operand_a_o[30]
port 90 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 alu_operand_a_o[31]
port 91 nsew signal output
rlabel metal3 s 199200 123768 200000 123888 6 alu_operand_a_o[32]
port 92 nsew signal output
rlabel metal2 s 160374 199200 160430 200000 6 alu_operand_a_o[3]
port 93 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 alu_operand_a_o[4]
port 94 nsew signal output
rlabel metal2 s 104990 199200 105046 200000 6 alu_operand_a_o[5]
port 95 nsew signal output
rlabel metal2 s 75366 199200 75422 200000 6 alu_operand_a_o[6]
port 96 nsew signal output
rlabel metal2 s 101770 199200 101826 200000 6 alu_operand_a_o[7]
port 97 nsew signal output
rlabel metal3 s 199200 47608 200000 47728 6 alu_operand_a_o[8]
port 98 nsew signal output
rlabel metal2 s 177118 199200 177174 200000 6 alu_operand_a_o[9]
port 99 nsew signal output
rlabel metal3 s 0 158448 800 158568 6 alu_operand_b_o[0]
port 100 nsew signal output
rlabel metal3 s 0 124448 800 124568 6 alu_operand_b_o[10]
port 101 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 alu_operand_b_o[11]
port 102 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 alu_operand_b_o[12]
port 103 nsew signal output
rlabel metal3 s 199200 74808 200000 74928 6 alu_operand_b_o[13]
port 104 nsew signal output
rlabel metal2 s 144274 199200 144330 200000 6 alu_operand_b_o[14]
port 105 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 alu_operand_b_o[15]
port 106 nsew signal output
rlabel metal3 s 0 68688 800 68808 6 alu_operand_b_o[16]
port 107 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 alu_operand_b_o[17]
port 108 nsew signal output
rlabel metal3 s 199200 175448 200000 175568 6 alu_operand_b_o[18]
port 109 nsew signal output
rlabel metal2 s 16762 199200 16818 200000 6 alu_operand_b_o[19]
port 110 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 alu_operand_b_o[1]
port 111 nsew signal output
rlabel metal2 s 199658 199200 199714 200000 6 alu_operand_b_o[20]
port 112 nsew signal output
rlabel metal3 s 199200 16328 200000 16448 6 alu_operand_b_o[21]
port 113 nsew signal output
rlabel metal3 s 0 189728 800 189848 6 alu_operand_b_o[22]
port 114 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 alu_operand_b_o[23]
port 115 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 alu_operand_b_o[24]
port 116 nsew signal output
rlabel metal3 s 0 127848 800 127968 6 alu_operand_b_o[25]
port 117 nsew signal output
rlabel metal2 s 114650 199200 114706 200000 6 alu_operand_b_o[26]
port 118 nsew signal output
rlabel metal3 s 199200 133968 200000 134088 6 alu_operand_b_o[27]
port 119 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 alu_operand_b_o[28]
port 120 nsew signal output
rlabel metal3 s 199200 189048 200000 189168 6 alu_operand_b_o[29]
port 121 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 alu_operand_b_o[2]
port 122 nsew signal output
rlabel metal2 s 46386 199200 46442 200000 6 alu_operand_b_o[30]
port 123 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 alu_operand_b_o[31]
port 124 nsew signal output
rlabel metal3 s 199200 33328 200000 33448 6 alu_operand_b_o[32]
port 125 nsew signal output
rlabel metal2 s 23202 199200 23258 200000 6 alu_operand_b_o[3]
port 126 nsew signal output
rlabel metal2 s 133970 0 134026 800 6 alu_operand_b_o[4]
port 127 nsew signal output
rlabel metal3 s 199200 192448 200000 192568 6 alu_operand_b_o[5]
port 128 nsew signal output
rlabel metal3 s 199200 109488 200000 109608 6 alu_operand_b_o[6]
port 129 nsew signal output
rlabel metal2 s 128174 199200 128230 200000 6 alu_operand_b_o[7]
port 130 nsew signal output
rlabel metal3 s 0 141448 800 141568 6 alu_operand_b_o[8]
port 131 nsew signal output
rlabel metal3 s 199200 195848 200000 195968 6 alu_operand_b_o[9]
port 132 nsew signal output
rlabel metal2 s 170034 0 170090 800 6 clk
port 133 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 div_en_i
port 134 nsew signal input
rlabel metal2 s 196438 0 196494 800 6 equal_to_zero
port 135 nsew signal input
rlabel metal3 s 199200 150968 200000 151088 6 mult_en_i
port 136 nsew signal input
rlabel metal3 s 0 179528 800 179648 6 multdiv_result_o[0]
port 137 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 multdiv_result_o[10]
port 138 nsew signal output
rlabel metal3 s 0 131248 800 131368 6 multdiv_result_o[11]
port 139 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 multdiv_result_o[12]
port 140 nsew signal output
rlabel metal3 s 199200 64608 200000 64728 6 multdiv_result_o[13]
port 141 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 multdiv_result_o[14]
port 142 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 multdiv_result_o[15]
port 143 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 multdiv_result_o[16]
port 144 nsew signal output
rlabel metal2 s 199658 0 199714 800 6 multdiv_result_o[17]
port 145 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 multdiv_result_o[18]
port 146 nsew signal output
rlabel metal3 s 199200 172048 200000 172168 6 multdiv_result_o[19]
port 147 nsew signal output
rlabel metal3 s 199200 127168 200000 127288 6 multdiv_result_o[1]
port 148 nsew signal output
rlabel metal3 s 0 148248 800 148368 6 multdiv_result_o[20]
port 149 nsew signal output
rlabel metal2 s 65706 199200 65762 200000 6 multdiv_result_o[21]
port 150 nsew signal output
rlabel metal2 s 192574 0 192630 800 6 multdiv_result_o[22]
port 151 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 multdiv_result_o[23]
port 152 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 multdiv_result_o[24]
port 153 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 multdiv_result_o[25]
port 154 nsew signal output
rlabel metal2 s 167458 199200 167514 200000 6 multdiv_result_o[26]
port 155 nsew signal output
rlabel metal3 s 199200 54408 200000 54528 6 multdiv_result_o[27]
port 156 nsew signal output
rlabel metal2 s 39302 199200 39358 200000 6 multdiv_result_o[28]
port 157 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 multdiv_result_o[29]
port 158 nsew signal output
rlabel metal2 s 10322 199200 10378 200000 6 multdiv_result_o[2]
port 159 nsew signal output
rlabel metal3 s 0 186328 800 186448 6 multdiv_result_o[30]
port 160 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 multdiv_result_o[31]
port 161 nsew signal output
rlabel metal3 s 199200 168648 200000 168768 6 multdiv_result_o[3]
port 162 nsew signal output
rlabel metal3 s 0 182928 800 183048 6 multdiv_result_o[4]
port 163 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 multdiv_result_o[5]
port 164 nsew signal output
rlabel metal2 s 26422 199200 26478 200000 6 multdiv_result_o[6]
port 165 nsew signal output
rlabel metal2 s 163594 0 163650 800 6 multdiv_result_o[7]
port 166 nsew signal output
rlabel metal3 s 199200 9528 200000 9648 6 multdiv_result_o[8]
port 167 nsew signal output
rlabel metal2 s 147494 199200 147550 200000 6 multdiv_result_o[9]
port 168 nsew signal output
rlabel metal3 s 199200 116288 200000 116408 6 op_a_i[0]
port 169 nsew signal input
rlabel metal2 s 52826 199200 52882 200000 6 op_a_i[10]
port 170 nsew signal input
rlabel metal2 s 62486 199200 62542 200000 6 op_a_i[11]
port 171 nsew signal input
rlabel metal2 s 56046 199200 56102 200000 6 op_a_i[12]
port 172 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 op_a_i[13]
port 173 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 op_a_i[14]
port 174 nsew signal input
rlabel metal3 s 0 144848 800 144968 6 op_a_i[15]
port 175 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 op_a_i[16]
port 176 nsew signal input
rlabel metal2 s 196438 199200 196494 200000 6 op_a_i[17]
port 177 nsew signal input
rlabel metal3 s 199200 161848 200000 161968 6 op_a_i[18]
port 178 nsew signal input
rlabel metal2 s 88890 199200 88946 200000 6 op_a_i[19]
port 179 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 op_a_i[1]
port 180 nsew signal input
rlabel metal3 s 199200 78888 200000 79008 6 op_a_i[20]
port 181 nsew signal input
rlabel metal3 s 0 120368 800 120488 6 op_a_i[21]
port 182 nsew signal input
rlabel metal2 s 3238 199200 3294 200000 6 op_a_i[22]
port 183 nsew signal input
rlabel metal3 s 199200 112888 200000 113008 6 op_a_i[23]
port 184 nsew signal input
rlabel metal3 s 0 161848 800 161968 6 op_a_i[24]
port 185 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 op_a_i[25]
port 186 nsew signal input
rlabel metal3 s 199200 185648 200000 185768 6 op_a_i[26]
port 187 nsew signal input
rlabel metal2 s 108210 199200 108266 200000 6 op_a_i[27]
port 188 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 op_a_i[28]
port 189 nsew signal input
rlabel metal3 s 199200 85688 200000 85808 6 op_a_i[29]
port 190 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 op_a_i[2]
port 191 nsew signal input
rlabel metal3 s 199200 29928 200000 30048 6 op_a_i[30]
port 192 nsew signal input
rlabel metal3 s 0 176128 800 176248 6 op_a_i[31]
port 193 nsew signal input
rlabel metal2 s 182914 0 182970 800 6 op_a_i[3]
port 194 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 op_a_i[4]
port 195 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 op_a_i[5]
port 196 nsew signal input
rlabel metal3 s 199200 57808 200000 57928 6 op_a_i[6]
port 197 nsew signal input
rlabel metal2 s 193218 199200 193274 200000 6 op_a_i[7]
port 198 nsew signal input
rlabel metal3 s 199200 147568 200000 147688 6 op_a_i[8]
port 199 nsew signal input
rlabel metal2 s 189354 0 189410 800 6 op_a_i[9]
port 200 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 op_b_i[0]
port 201 nsew signal input
rlabel metal3 s 199200 89088 200000 89208 6 op_b_i[10]
port 202 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 op_b_i[11]
port 203 nsew signal input
rlabel metal3 s 199200 157768 200000 157888 6 op_b_i[12]
port 204 nsew signal input
rlabel metal2 s 180338 199200 180394 200000 6 op_b_i[13]
port 205 nsew signal input
rlabel metal3 s 199200 2728 200000 2848 6 op_b_i[14]
port 206 nsew signal input
rlabel metal2 s 173898 199200 173954 200000 6 op_b_i[15]
port 207 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 op_b_i[16]
port 208 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 op_b_i[17]
port 209 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 op_b_i[18]
port 210 nsew signal input
rlabel metal2 s 18 0 74 800 6 op_b_i[19]
port 211 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 op_b_i[1]
port 212 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 op_b_i[20]
port 213 nsew signal input
rlabel metal2 s 7102 199200 7158 200000 6 op_b_i[21]
port 214 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 op_b_i[22]
port 215 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 op_b_i[23]
port 216 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 op_b_i[24]
port 217 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 op_b_i[25]
port 218 nsew signal input
rlabel metal2 s 124954 199200 125010 200000 6 op_b_i[26]
port 219 nsew signal input
rlabel metal2 s 81806 199200 81862 200000 6 op_b_i[27]
port 220 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 op_b_i[28]
port 221 nsew signal input
rlabel metal2 s 153934 199200 153990 200000 6 op_b_i[29]
port 222 nsew signal input
rlabel metal3 s 199200 44208 200000 44328 6 op_b_i[2]
port 223 nsew signal input
rlabel metal3 s 0 151648 800 151768 6 op_b_i[30]
port 224 nsew signal input
rlabel metal3 s 199200 144168 200000 144288 6 op_b_i[31]
port 225 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 op_b_i[3]
port 226 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 op_b_i[4]
port 227 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 op_b_i[5]
port 228 nsew signal input
rlabel metal3 s 199200 140768 200000 140888 6 op_b_i[6]
port 229 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 op_b_i[7]
port 230 nsew signal input
rlabel metal2 s 141054 199200 141110 200000 6 op_b_i[8]
port 231 nsew signal input
rlabel metal2 s 137834 199200 137890 200000 6 op_b_i[9]
port 232 nsew signal input
rlabel metal3 s 0 196528 800 196648 6 operator_i[0]
port 233 nsew signal input
rlabel metal2 s 29642 199200 29698 200000 6 operator_i[1]
port 234 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 ready_o
port 235 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 rst_n
port 236 nsew signal input
rlabel metal3 s 0 172728 800 172848 6 signed_mode_i[0]
port 237 nsew signal input
rlabel metal3 s 199200 95888 200000 96008 6 signed_mode_i[1]
port 238 nsew signal input
rlabel metal5 s 1104 5298 198812 5618 6 vccd1
port 239 nsew power input
rlabel metal5 s 1104 35934 198812 36254 6 vccd1
port 239 nsew power input
rlabel metal5 s 1104 66570 198812 66890 6 vccd1
port 239 nsew power input
rlabel metal5 s 1104 97206 198812 97526 6 vccd1
port 239 nsew power input
rlabel metal5 s 1104 127842 198812 128162 6 vccd1
port 239 nsew power input
rlabel metal5 s 1104 158478 198812 158798 6 vccd1
port 239 nsew power input
rlabel metal5 s 1104 189114 198812 189434 6 vccd1
port 239 nsew power input
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 239 nsew power input
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 239 nsew power input
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 239 nsew power input
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 239 nsew power input
rlabel metal4 s 127088 2128 127408 197520 6 vccd1
port 239 nsew power input
rlabel metal4 s 157808 2128 158128 197520 6 vccd1
port 239 nsew power input
rlabel metal4 s 188528 2128 188848 197520 6 vccd1
port 239 nsew power input
rlabel metal5 s 1104 20616 198812 20936 6 vssd1
port 240 nsew ground input
rlabel metal5 s 1104 51252 198812 51572 6 vssd1
port 240 nsew ground input
rlabel metal5 s 1104 81888 198812 82208 6 vssd1
port 240 nsew ground input
rlabel metal5 s 1104 112524 198812 112844 6 vssd1
port 240 nsew ground input
rlabel metal5 s 1104 143160 198812 143480 6 vssd1
port 240 nsew ground input
rlabel metal5 s 1104 173796 198812 174116 6 vssd1
port 240 nsew ground input
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 240 nsew ground input
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 240 nsew ground input
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 240 nsew ground input
rlabel metal4 s 111728 2128 112048 197520 6 vssd1
port 240 nsew ground input
rlabel metal4 s 142448 2128 142768 197520 6 vssd1
port 240 nsew ground input
rlabel metal4 s 173168 2128 173488 197520 6 vssd1
port 240 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 200000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 21152680
string GDS_FILE /home/mbaykenar/Desktop/first_asic/openlane/zeroriscy_multdiv_fast/runs/zeroriscy_multdiv_fast/results/finishing/zeroriscy_multdiv_fast.magic.gds
string GDS_START 1106636
<< end >>

